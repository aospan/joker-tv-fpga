
module probe (
	probe,
	source);	

	input	[510:0]	probe;
	output	[31:0]	source;
endmodule
