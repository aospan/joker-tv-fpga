parameter	[7:0]	DESCR_USB2_DEVICE	= 'd0;
parameter	[6:0]	DESCR_USB3_DEVICE	= 'd0;
parameter	[7:0]	DESCR_USB2_DEVICE_QUAL	= 'd18;
parameter	[7:0]	DESCR_USB2_CONFIG	= 'd28;
parameter	[6:0]	DESCR_USB3_CONFIG	= 'd5;
parameter	[7:0]	DESCR_USB2_CONFIG_LEN	= 'd48;
parameter	[6:0]	DESCR_USB3_CONFIG_LEN	= 'd66;
parameter	[6:0]	DESCR_USB3_BOS    	= 'd22;
parameter	[6:0]	DESCR_USB3_BOS_LEN	= 'd22;
parameter	[7:0]	DESCR_USB2_STRING0	= 'd76;
parameter	[6:0]	DESCR_USB3_STRING0	= 'd28;
parameter	[7:0]	DESCR_USB2_STRING1	= 'd80;
parameter	[6:0]	DESCR_USB3_STRING1	= 'd29;
parameter	[7:0]	DESCR_USB2_STRING2	= 'd118;
parameter	[6:0]	DESCR_USB3_STRING2	= 'd39;
parameter	[7:0]	DESCR_USB2_STRING3	= 'd136;
parameter	[6:0]	DESCR_USB3_STRING3	= 'd44;
parameter	[7:0]	DESCR_USB2_CONFUNSET	= 'd158;
parameter	[6:0]	DESCR_USB3_CONFUNSET	= 'd50;
parameter	[7:0]	DESCR_USB2_CONFSET	= 'd159;
parameter	[6:0]	DESCR_USB3_CONFSET	= 'd51;
parameter	[7:0]	DESCR_USB2_EOF     	= 'd160;
parameter	[6:0]	DESCR_USB3_EOF     	= 'd52;
