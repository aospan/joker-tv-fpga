parameter	[7:0]	DESCR_USB2_DEVICE	= 'd0;
parameter	[6:0]	DESCR_USB3_DEVICE	= 'd0;
parameter	[7:0]	DESCR_USB2_DEVICE_QUAL	= 'd18;
parameter	[7:0]	DESCR_USB2_CONFIG	= 'd28;
parameter	[6:0]	DESCR_USB3_CONFIG	= 'd5;
parameter	[7:0]	DESCR_USB2_CONFIG_LEN	= 'd48;
parameter	[6:0]	DESCR_USB3_CONFIG_LEN	= 'd66;
parameter	[6:0]	DESCR_USB3_BOS    	= 'd22;
parameter	[6:0]	DESCR_USB3_BOS_LEN	= 'd22;
parameter	[7:0]	DESCR_USB2_STRING0	= 'd76;
parameter	[6:0]	DESCR_USB3_STRING0	= 'd28;
parameter	[7:0]	DESCR_USB2_STRING1	= 'd82;
parameter	[6:0]	DESCR_USB3_STRING1	= 'd30;
parameter	[7:0]	DESCR_USB2_STRING2	= 'd120;
parameter	[6:0]	DESCR_USB3_STRING2	= 'd40;
parameter	[7:0]	DESCR_USB2_STRING3	= 'd138;
parameter	[6:0]	DESCR_USB3_STRING3	= 'd45;
parameter	[7:0]	DESCR_USB2_STRING238	= 'd160;
parameter	[6:0]	DESCR_USB3_STRING238	= 'd51;
parameter	[7:0]	DESCR_USB2_MS_COMPAT	= 'd178;
parameter	[6:0]	DESCR_USB3_MS_COMPAT	= 'd56;
parameter	[7:0]	DESCR_USB2_CONFUNSET	= 'd218;
parameter	[6:0]	DESCR_USB3_CONFUNSET	= 'd66;
parameter	[7:0]	DESCR_USB2_CONFSET	= 'd219;
parameter	[6:0]	DESCR_USB3_CONFSET	= 'd67;
parameter	[7:0]	DESCR_USB2_STATUS	= 'd220;
parameter	[6:0]	DESCR_USB3_STATUS	= 'd68;
parameter	[7:0]	DESCR_USB2_EOF     	= 'd222;
parameter	[6:0]	DESCR_USB3_EOF     	= 'd69;
