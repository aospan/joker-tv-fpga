parameter	[7:0]	DESCR_USB2_DEVICE	= 'd0;
parameter	[6:0]	DESCR_USB3_DEVICE	= 'd0;
parameter	[7:0]	DESCR_USB2_DEVICE_QUAL	= 'd18;
parameter	[7:0]	DESCR_USB2_CONFIG	= 'd28;
parameter	[6:0]	DESCR_USB3_CONFIG	= 'd5;
parameter	[7:0]	DESCR_USB2_CONFIG_LEN	= 'd55;
parameter	[6:0]	DESCR_USB3_CONFIG_LEN	= 'd79;
parameter	[6:0]	DESCR_USB3_BOS    	= 'd25;
parameter	[6:0]	DESCR_USB3_BOS_LEN	= 'd22;
parameter	[7:0]	DESCR_USB2_STRING0	= 'd83;
parameter	[6:0]	DESCR_USB3_STRING0	= 'd31;
parameter	[7:0]	DESCR_USB2_STRING1	= 'd89;
parameter	[6:0]	DESCR_USB3_STRING1	= 'd33;
parameter	[7:0]	DESCR_USB2_STRING2	= 'd127;
parameter	[6:0]	DESCR_USB3_STRING2	= 'd43;
parameter	[7:0]	DESCR_USB2_STRING3	= 'd145;
parameter	[6:0]	DESCR_USB3_STRING3	= 'd48;
parameter	[7:0]	DESCR_USB2_STRING238	= 'd167;
parameter	[6:0]	DESCR_USB3_STRING238	= 'd54;
parameter	[7:0]	DESCR_USB2_MS_COMPAT	= 'd185;
parameter	[6:0]	DESCR_USB3_MS_COMPAT	= 'd59;
parameter	[7:0]	DESCR_USB2_CONFUNSET	= 'd225;
parameter	[6:0]	DESCR_USB3_CONFUNSET	= 'd69;
parameter	[7:0]	DESCR_USB2_CONFSET	= 'd226;
parameter	[6:0]	DESCR_USB3_CONFSET	= 'd70;
parameter	[7:0]	DESCR_USB2_STATUS	= 'd227;
parameter	[6:0]	DESCR_USB3_STATUS	= 'd71;
parameter	[7:0]	DESCR_USB2_EOF     	= 'd229;
parameter	[6:0]	DESCR_USB3_EOF     	= 'd72;
